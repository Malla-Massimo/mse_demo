// base_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module base_system (
		input  wire [9:0]  cam_data,      //       cam.data
		input  wire        cam_hsync,     //          .hsync
		input  wire        cam_pxlclk,    //          .pxlclk
		output wire        cam_pwrdwn,    //          .pwrdwn
		output wire        cam_rstb,      //          .rstb
		input  wire        cam_vsync,     //          .vsync
		input  wire        clk_clk,       //       clk.clk
		output wire        dac_clk_clk,   //   dac_clk.clk
		input  wire [7:0]  dipsw_export,  //     dipsw.export
		output wire        i2c_scl,       //       i2c.scl
		inout  wire        i2c_sda,       //          .sda
		output wire        lcd_csb,       //       lcd.csb
		inout  wire [15:0] lcd_db,        //          .db
		output wire        lcd_dcb,       //          .dcb
		output wire        lcd_im,        //          .im
		output wire        lcd_rb,        //          .rb
		output wire        lcd_resb,      //          .resb
		output wire        lcd_wb,        //          .wb
		output wire        mclk_clk,      //      mclk.clk
		input  wire        reset_reset_n, //     reset.reset_n
		output wire [11:0] sdram_addr,    //     sdram.addr
		output wire [1:0]  sdram_ba,      //          .ba
		output wire        sdram_cas_n,   //          .cas_n
		output wire        sdram_cke,     //          .cke
		output wire        sdram_cs_n,    //          .cs_n
		inout  wire [15:0] sdram_dq,      //          .dq
		output wire [1:0]  sdram_dqm,     //          .dqm
		output wire        sdram_ras_n,   //          .ras_n
		output wire        sdram_we_n,    //          .we_n
		output wire        sdram_clk_clk, // sdram_clk.clk
		output wire [9:0]  vga_blue,      //       vga.blue
		output wire [9:0]  vga_green,     //          .green
		output wire        vga_hsync,     //          .hsync
		output wire [9:0]  vga_red,       //          .red
		output wire        vga_vsync      //          .vsync
	);

	wire         altpll_0_c0_clk;                                            // altpll_0:c0 -> [ProfileTimer:clk, Systimer:clk, cam_ctrl:Clock, i2c_ctrl:clock, irq_mapper:clk, jtag_uart:clk, lcd_ctrl:Clock, mm_interconnect_0:altpll_0_c0_clk, nios2_gen2_0:clk, pio_0:clk, rst_controller:clk, sdram_ctrl:clk, sysid:clock, vga_dma_0:Clock]
	wire         altpll_0_c4_clk;                                            // altpll_0:c4 -> vga_dma_0:PixelClock
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [24:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                     // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire   [3:0] nios2_gen2_0_data_master_burstcount;                        // nios2_gen2_0:d_burstcount -> mm_interconnect_0:nios2_gen2_0_data_master_burstcount
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [24:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;              // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire   [3:0] nios2_gen2_0_instruction_master_burstcount;                 // nios2_gen2_0:i_burstcount -> mm_interconnect_0:nios2_gen2_0_instruction_master_burstcount
	wire  [31:0] lcd_ctrl_master_readdata;                                   // mm_interconnect_0:lcd_ctrl_master_readdata -> lcd_ctrl:master_read_data
	wire         lcd_ctrl_master_waitrequest;                                // mm_interconnect_0:lcd_ctrl_master_waitrequest -> lcd_ctrl:master_wait_request
	wire  [31:0] lcd_ctrl_master_address;                                    // lcd_ctrl:master_address -> mm_interconnect_0:lcd_ctrl_master_address
	wire         lcd_ctrl_master_read;                                       // lcd_ctrl:master_read -> mm_interconnect_0:lcd_ctrl_master_read
	wire         lcd_ctrl_master_readdatavalid;                              // mm_interconnect_0:lcd_ctrl_master_readdatavalid -> lcd_ctrl:master_read_data_valid
	wire   [7:0] lcd_ctrl_master_burstcount;                                 // lcd_ctrl:master_burst_count -> mm_interconnect_0:lcd_ctrl_master_burstcount
	wire         cam_ctrl_master_waitrequest;                                // mm_interconnect_0:cam_ctrl_master_waitrequest -> cam_ctrl:master_wait_req
	wire  [31:0] cam_ctrl_master_address;                                    // cam_ctrl:master_address -> mm_interconnect_0:cam_ctrl_master_address
	wire         cam_ctrl_master_write;                                      // cam_ctrl:master_we -> mm_interconnect_0:cam_ctrl_master_write
	wire  [31:0] cam_ctrl_master_writedata;                                  // cam_ctrl:master_write_data -> mm_interconnect_0:cam_ctrl_master_writedata
	wire   [9:0] cam_ctrl_master_burstcount;                                 // cam_ctrl:master_burst_count -> mm_interconnect_0:cam_ctrl_master_burstcount
	wire  [31:0] vga_dma_0_master_readdata;                                  // mm_interconnect_0:vga_dma_0_master_readdata -> vga_dma_0:master_read_data
	wire         vga_dma_0_master_waitrequest;                               // mm_interconnect_0:vga_dma_0_master_waitrequest -> vga_dma_0:master_waitrequest
	wire  [31:0] vga_dma_0_master_address;                                   // vga_dma_0:master_address -> mm_interconnect_0:vga_dma_0_master_address
	wire         vga_dma_0_master_read;                                      // vga_dma_0:master_read -> mm_interconnect_0:vga_dma_0_master_read
	wire         vga_dma_0_master_readdatavalid;                             // mm_interconnect_0:vga_dma_0_master_readdatavalid -> vga_dma_0:master_data_valid
	wire   [9:0] vga_dma_0_master_burstcount;                                // vga_dma_0:master_burstcount -> mm_interconnect_0:vga_dma_0_master_burstcount
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;             // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;              // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;              // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;               // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                  // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                 // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;             // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_sdram_ctrl_s1_chipselect;                 // mm_interconnect_0:sdram_ctrl_s1_chipselect -> sdram_ctrl:az_cs
	wire  [15:0] mm_interconnect_0_sdram_ctrl_s1_readdata;                   // sdram_ctrl:za_data -> mm_interconnect_0:sdram_ctrl_s1_readdata
	wire         mm_interconnect_0_sdram_ctrl_s1_waitrequest;                // sdram_ctrl:za_waitrequest -> mm_interconnect_0:sdram_ctrl_s1_waitrequest
	wire  [22:0] mm_interconnect_0_sdram_ctrl_s1_address;                    // mm_interconnect_0:sdram_ctrl_s1_address -> sdram_ctrl:az_addr
	wire         mm_interconnect_0_sdram_ctrl_s1_read;                       // mm_interconnect_0:sdram_ctrl_s1_read -> sdram_ctrl:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_ctrl_s1_byteenable;                 // mm_interconnect_0:sdram_ctrl_s1_byteenable -> sdram_ctrl:az_be_n
	wire         mm_interconnect_0_sdram_ctrl_s1_readdatavalid;              // sdram_ctrl:za_valid -> mm_interconnect_0:sdram_ctrl_s1_readdatavalid
	wire         mm_interconnect_0_sdram_ctrl_s1_write;                      // mm_interconnect_0:sdram_ctrl_s1_write -> sdram_ctrl:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_ctrl_s1_writedata;                  // mm_interconnect_0:sdram_ctrl_s1_writedata -> sdram_ctrl:az_data
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                        // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                         // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_systimer_s1_chipselect;                   // mm_interconnect_0:Systimer_s1_chipselect -> Systimer:chipselect
	wire  [15:0] mm_interconnect_0_systimer_s1_readdata;                     // Systimer:readdata -> mm_interconnect_0:Systimer_s1_readdata
	wire   [2:0] mm_interconnect_0_systimer_s1_address;                      // mm_interconnect_0:Systimer_s1_address -> Systimer:address
	wire         mm_interconnect_0_systimer_s1_write;                        // mm_interconnect_0:Systimer_s1_write -> Systimer:write_n
	wire  [15:0] mm_interconnect_0_systimer_s1_writedata;                    // mm_interconnect_0:Systimer_s1_writedata -> Systimer:writedata
	wire         mm_interconnect_0_profiletimer_s1_chipselect;               // mm_interconnect_0:ProfileTimer_s1_chipselect -> ProfileTimer:chipselect
	wire  [15:0] mm_interconnect_0_profiletimer_s1_readdata;                 // ProfileTimer:readdata -> mm_interconnect_0:ProfileTimer_s1_readdata
	wire   [2:0] mm_interconnect_0_profiletimer_s1_address;                  // mm_interconnect_0:ProfileTimer_s1_address -> ProfileTimer:address
	wire         mm_interconnect_0_profiletimer_s1_write;                    // mm_interconnect_0:ProfileTimer_s1_write -> ProfileTimer:write_n
	wire  [15:0] mm_interconnect_0_profiletimer_s1_writedata;                // mm_interconnect_0:ProfileTimer_s1_writedata -> ProfileTimer:writedata
	wire         mm_interconnect_0_lcd_ctrl_slave_chipselect;                // mm_interconnect_0:lcd_ctrl_slave_chipselect -> lcd_ctrl:slave_cs
	wire  [31:0] mm_interconnect_0_lcd_ctrl_slave_readdata;                  // lcd_ctrl:slave_read_data -> mm_interconnect_0:lcd_ctrl_slave_readdata
	wire         mm_interconnect_0_lcd_ctrl_slave_waitrequest;               // lcd_ctrl:slave_wait_request -> mm_interconnect_0:lcd_ctrl_slave_waitrequest
	wire   [2:0] mm_interconnect_0_lcd_ctrl_slave_address;                   // mm_interconnect_0:lcd_ctrl_slave_address -> lcd_ctrl:slave_address
	wire         mm_interconnect_0_lcd_ctrl_slave_read;                      // mm_interconnect_0:lcd_ctrl_slave_read -> lcd_ctrl:slave_rd
	wire         mm_interconnect_0_lcd_ctrl_slave_write;                     // mm_interconnect_0:lcd_ctrl_slave_write -> lcd_ctrl:slave_we
	wire  [31:0] mm_interconnect_0_lcd_ctrl_slave_writedata;                 // mm_interconnect_0:lcd_ctrl_slave_writedata -> lcd_ctrl:slave_write_data
	wire         mm_interconnect_0_i2c_ctrl_slave_chipselect;                // mm_interconnect_0:i2c_ctrl_slave_chipselect -> i2c_ctrl:slave_cs
	wire  [31:0] mm_interconnect_0_i2c_ctrl_slave_readdata;                  // i2c_ctrl:slave_read_data -> mm_interconnect_0:i2c_ctrl_slave_readdata
	wire   [1:0] mm_interconnect_0_i2c_ctrl_slave_address;                   // mm_interconnect_0:i2c_ctrl_slave_address -> i2c_ctrl:slave_address
	wire   [3:0] mm_interconnect_0_i2c_ctrl_slave_byteenable;                // mm_interconnect_0:i2c_ctrl_slave_byteenable -> i2c_ctrl:slave_byte_enables
	wire         mm_interconnect_0_i2c_ctrl_slave_write;                     // mm_interconnect_0:i2c_ctrl_slave_write -> i2c_ctrl:slave_we
	wire  [31:0] mm_interconnect_0_i2c_ctrl_slave_writedata;                 // mm_interconnect_0:i2c_ctrl_slave_writedata -> i2c_ctrl:slave_write_data
	wire         mm_interconnect_0_cam_ctrl_slave_chipselect;                // mm_interconnect_0:cam_ctrl_slave_chipselect -> cam_ctrl:slave_cs
	wire  [31:0] mm_interconnect_0_cam_ctrl_slave_readdata;                  // cam_ctrl:slave_read_data -> mm_interconnect_0:cam_ctrl_slave_readdata
	wire   [2:0] mm_interconnect_0_cam_ctrl_slave_address;                   // mm_interconnect_0:cam_ctrl_slave_address -> cam_ctrl:slave_address
	wire         mm_interconnect_0_cam_ctrl_slave_write;                     // mm_interconnect_0:cam_ctrl_slave_write -> cam_ctrl:slave_we
	wire  [31:0] mm_interconnect_0_cam_ctrl_slave_writedata;                 // mm_interconnect_0:cam_ctrl_slave_writedata -> cam_ctrl:slave_write_data
	wire         mm_interconnect_0_vga_dma_0_slave_chipselect;               // mm_interconnect_0:vga_dma_0_slave_chipselect -> vga_dma_0:slave_cs
	wire   [0:0] mm_interconnect_0_vga_dma_0_slave_address;                  // mm_interconnect_0:vga_dma_0_slave_address -> vga_dma_0:slave_address
	wire         mm_interconnect_0_vga_dma_0_slave_write;                    // mm_interconnect_0:vga_dma_0_slave_write -> vga_dma_0:slave_we
	wire  [31:0] mm_interconnect_0_vga_dma_0_slave_writedata;                // mm_interconnect_0:vga_dma_0_slave_writedata -> vga_dma_0:slave_write_data
	wire         irq_mapper_receiver0_irq;                                   // cam_ctrl:IRQ -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // lcd_ctrl:end_of_transaction_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                   // i2c_ctrl:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                   // Systimer:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                   // ProfileTimer:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [ProfileTimer:reset_n, Systimer:reset_n, cam_ctrl:Reset, i2c_ctrl:reset, irq_mapper:reset, jtag_uart:rst_n, lcd_ctrl:Reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, pio_0:reset_n, rst_translator:in_reset, sdram_ctrl:reset_n, sysid:reset_n, vga_dma_0:Reset]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]

	base_system_ProfileTimer profiletimer (
		.clk        (altpll_0_c0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_profiletimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_profiletimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_profiletimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_profiletimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_profiletimer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                      //   irq.irq
	);

	base_system_ProfileTimer systimer (
		.clk        (altpll_0_c0_clk),                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_systimer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                  //   irq.irq
	);

	base_system_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (mclk_clk),                                       //                    c1.clk
		.c2                 (sdram_clk_clk),                                  //                    c2.clk
		.c3                 (dac_clk_clk),                                    //                    c3.clk
		.c4                 (altpll_0_c4_clk),                                //                    c4.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0),                                           //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          ()                                                //           (terminated)
	);

	cam_dma cam_ctrl (
		.Reset              (rst_controller_reset_out_reset),              //     reset.reset
		.slave_address      (mm_interconnect_0_cam_ctrl_slave_address),    //     slave.address
		.slave_cs           (mm_interconnect_0_cam_ctrl_slave_chipselect), //          .chipselect
		.slave_read_data    (mm_interconnect_0_cam_ctrl_slave_readdata),   //          .readdata
		.slave_we           (mm_interconnect_0_cam_ctrl_slave_write),      //          .write
		.slave_write_data   (mm_interconnect_0_cam_ctrl_slave_writedata),  //          .writedata
		.Clock              (altpll_0_c0_clk),                             //     clock.clk
		.IRQ                (irq_mapper_receiver0_irq),                    // interrupt.irq
		.DataIn             (cam_data),                                    //    camera.data
		.HSync              (cam_hsync),                                   //          .hsync
		.PixelClk           (cam_pxlclk),                                  //          .pxlclk
		.PowerDown          (cam_pwrdwn),                                  //          .pwrdwn
		.ResetBar           (cam_rstb),                                    //          .rstb
		.VSync              (cam_vsync),                                   //          .vsync
		.master_address     (cam_ctrl_master_address),                     //    master.address
		.master_burst_count (cam_ctrl_master_burstcount),                  //          .burstcount
		.master_wait_req    (cam_ctrl_master_waitrequest),                 //          .waitrequest
		.master_we          (cam_ctrl_master_write),                       //          .write
		.master_write_data  (cam_ctrl_master_writedata)                    //          .writedata
	);

	i2c_core i2c_ctrl (
		.reset              (rst_controller_reset_out_reset),              //    reset.reset
		.slave_address      (mm_interconnect_0_i2c_ctrl_slave_address),    //    slave.address
		.slave_byte_enables (mm_interconnect_0_i2c_ctrl_slave_byteenable), //         .byteenable
		.slave_cs           (mm_interconnect_0_i2c_ctrl_slave_chipselect), //         .chipselect
		.slave_read_data    (mm_interconnect_0_i2c_ctrl_slave_readdata),   //         .readdata
		.slave_we           (mm_interconnect_0_i2c_ctrl_slave_write),      //         .write
		.slave_write_data   (mm_interconnect_0_i2c_ctrl_slave_writedata),  //         .writedata
		.clock              (altpll_0_c0_clk),                             //    clock.clk
		.SCL                (i2c_scl),                                     // i2c_port.scl
		.SDA                (i2c_sda),                                     //         .sda
		.irq                (irq_mapper_receiver3_irq)                     //      irq.irq
	);

	base_system_jtag_uart jtag_uart (
		.clk            (altpll_0_c0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	lcd_dma lcd_ctrl (
		.Reset                  (rst_controller_reset_out_reset),               //    reset.reset
		.slave_address          (mm_interconnect_0_lcd_ctrl_slave_address),     //    slave.address
		.slave_cs               (mm_interconnect_0_lcd_ctrl_slave_chipselect),  //         .chipselect
		.slave_rd               (mm_interconnect_0_lcd_ctrl_slave_read),        //         .read
		.slave_read_data        (mm_interconnect_0_lcd_ctrl_slave_readdata),    //         .readdata
		.slave_wait_request     (mm_interconnect_0_lcd_ctrl_slave_waitrequest), //         .waitrequest
		.slave_we               (mm_interconnect_0_lcd_ctrl_slave_write),       //         .write
		.slave_write_data       (mm_interconnect_0_lcd_ctrl_slave_writedata),   //         .writedata
		.master_read_data_valid (lcd_ctrl_master_readdatavalid),                //   master.readdatavalid
		.master_address         (lcd_ctrl_master_address),                      //         .address
		.master_burst_count     (lcd_ctrl_master_burstcount),                   //         .burstcount
		.master_read            (lcd_ctrl_master_read),                         //         .read
		.master_read_data       (lcd_ctrl_master_readdata),                     //         .readdata
		.master_wait_request    (lcd_ctrl_master_waitrequest),                  //         .waitrequest
		.Clock                  (altpll_0_c0_clk),                              //    clock.clk
		.ChipSelectBar          (lcd_csb),                                      // external.csb
		.DataBus                (lcd_db),                                       //         .db
		.DataCommandBar         (lcd_dcb),                                      //         .dcb
		.IM0                    (lcd_im),                                       //         .im
		.ReadBar                (lcd_rb),                                       //         .rb
		.ResetBar               (lcd_resb),                                     //         .resb
		.WriteBar               (lcd_wb),                                       //         .wb
		.end_of_transaction_irq (irq_mapper_receiver2_irq)                      //      irq.irq
	);

	base_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_burstcount                        (nios2_gen2_0_data_master_burstcount),                        //                          .burstcount
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_burstcount                        (nios2_gen2_0_instruction_master_burstcount),                 //                          .burstcount
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	base_system_pio_0 pio_0 (
		.clk      (altpll_0_c0_clk),                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_0_s1_readdata), //                    .readdata
		.in_port  (dipsw_export)                         // external_connection.export
	);

	base_system_sdram_ctrl sdram_ctrl (
		.clk            (altpll_0_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),               // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_ctrl_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_ctrl_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_ctrl_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_ctrl_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_ctrl_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_ctrl_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_ctrl_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_ctrl_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_ctrl_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                    //  wire.export
		.zs_ba          (sdram_ba),                                      //      .export
		.zs_cas_n       (sdram_cas_n),                                   //      .export
		.zs_cke         (sdram_cke),                                     //      .export
		.zs_cs_n        (sdram_cs_n),                                    //      .export
		.zs_dq          (sdram_dq),                                      //      .export
		.zs_dqm         (sdram_dqm),                                     //      .export
		.zs_ras_n       (sdram_ras_n),                                   //      .export
		.zs_we_n        (sdram_we_n)                                     //      .export
	);

	base_system_sysid sysid (
		.clock    (altpll_0_c0_clk),                                //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	vga_dma vga_dma_0 (
		.Reset              (rst_controller_reset_out_reset),               //    reset.reset
		.slave_address      (mm_interconnect_0_vga_dma_0_slave_address),    //    slave.address
		.slave_cs           (mm_interconnect_0_vga_dma_0_slave_chipselect), //         .chipselect
		.slave_we           (mm_interconnect_0_vga_dma_0_slave_write),      //         .write
		.slave_write_data   (mm_interconnect_0_vga_dma_0_slave_writedata),  //         .writedata
		.Clock              (altpll_0_c0_clk),                              //    clock.clk
		.PixelClock         (altpll_0_c4_clk),                              // pixelclk.clk
		.master_address     (vga_dma_0_master_address),                     //   master.address
		.master_burstcount  (vga_dma_0_master_burstcount),                  //         .burstcount
		.master_data_valid  (vga_dma_0_master_readdatavalid),               //         .readdatavalid
		.master_read        (vga_dma_0_master_read),                        //         .read
		.master_read_data   (vga_dma_0_master_readdata),                    //         .readdata
		.master_waitrequest (vga_dma_0_master_waitrequest),                 //         .waitrequest
		.blue               (vga_blue),                                     //      vga.blue
		.green              (vga_green),                                    //         .green
		.hsync              (vga_hsync),                                    //         .hsync
		.red                (vga_red),                                      //         .red
		.vsync              (vga_vsync)                                     //         .vsync
	);

	base_system_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                            //                                          altpll_0_c0.clk
		.clk_0_clk_clk                                              (clk_clk),                                                    //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                             //             nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.cam_ctrl_master_address                                    (cam_ctrl_master_address),                                    //                                      cam_ctrl_master.address
		.cam_ctrl_master_waitrequest                                (cam_ctrl_master_waitrequest),                                //                                                     .waitrequest
		.cam_ctrl_master_burstcount                                 (cam_ctrl_master_burstcount),                                 //                                                     .burstcount
		.cam_ctrl_master_write                                      (cam_ctrl_master_write),                                      //                                                     .write
		.cam_ctrl_master_writedata                                  (cam_ctrl_master_writedata),                                  //                                                     .writedata
		.lcd_ctrl_master_address                                    (lcd_ctrl_master_address),                                    //                                      lcd_ctrl_master.address
		.lcd_ctrl_master_waitrequest                                (lcd_ctrl_master_waitrequest),                                //                                                     .waitrequest
		.lcd_ctrl_master_burstcount                                 (lcd_ctrl_master_burstcount),                                 //                                                     .burstcount
		.lcd_ctrl_master_read                                       (lcd_ctrl_master_read),                                       //                                                     .read
		.lcd_ctrl_master_readdata                                   (lcd_ctrl_master_readdata),                                   //                                                     .readdata
		.lcd_ctrl_master_readdatavalid                              (lcd_ctrl_master_readdatavalid),                              //                                                     .readdatavalid
		.nios2_gen2_0_data_master_address                           (nios2_gen2_0_data_master_address),                           //                             nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                                                     .waitrequest
		.nios2_gen2_0_data_master_burstcount                        (nios2_gen2_0_data_master_burstcount),                        //                                                     .burstcount
		.nios2_gen2_0_data_master_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                                                     .byteenable
		.nios2_gen2_0_data_master_read                              (nios2_gen2_0_data_master_read),                              //                                                     .read
		.nios2_gen2_0_data_master_readdata                          (nios2_gen2_0_data_master_readdata),                          //                                                     .readdata
		.nios2_gen2_0_data_master_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                                                     .readdatavalid
		.nios2_gen2_0_data_master_write                             (nios2_gen2_0_data_master_write),                             //                                                     .write
		.nios2_gen2_0_data_master_writedata                         (nios2_gen2_0_data_master_writedata),                         //                                                     .writedata
		.nios2_gen2_0_data_master_debugaccess                       (nios2_gen2_0_data_master_debugaccess),                       //                                                     .debugaccess
		.nios2_gen2_0_instruction_master_address                    (nios2_gen2_0_instruction_master_address),                    //                      nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                (nios2_gen2_0_instruction_master_waitrequest),                //                                                     .waitrequest
		.nios2_gen2_0_instruction_master_burstcount                 (nios2_gen2_0_instruction_master_burstcount),                 //                                                     .burstcount
		.nios2_gen2_0_instruction_master_read                       (nios2_gen2_0_instruction_master_read),                       //                                                     .read
		.nios2_gen2_0_instruction_master_readdata                   (nios2_gen2_0_instruction_master_readdata),                   //                                                     .readdata
		.nios2_gen2_0_instruction_master_readdatavalid              (nios2_gen2_0_instruction_master_readdatavalid),              //                                                     .readdatavalid
		.vga_dma_0_master_address                                   (vga_dma_0_master_address),                                   //                                     vga_dma_0_master.address
		.vga_dma_0_master_waitrequest                               (vga_dma_0_master_waitrequest),                               //                                                     .waitrequest
		.vga_dma_0_master_burstcount                                (vga_dma_0_master_burstcount),                                //                                                     .burstcount
		.vga_dma_0_master_read                                      (vga_dma_0_master_read),                                      //                                                     .read
		.vga_dma_0_master_readdata                                  (vga_dma_0_master_readdata),                                  //                                                     .readdata
		.vga_dma_0_master_readdatavalid                             (vga_dma_0_master_readdatavalid),                             //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),               //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                 //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                  //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),              //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),             //                                                     .writedata
		.cam_ctrl_slave_address                                     (mm_interconnect_0_cam_ctrl_slave_address),                   //                                       cam_ctrl_slave.address
		.cam_ctrl_slave_write                                       (mm_interconnect_0_cam_ctrl_slave_write),                     //                                                     .write
		.cam_ctrl_slave_readdata                                    (mm_interconnect_0_cam_ctrl_slave_readdata),                  //                                                     .readdata
		.cam_ctrl_slave_writedata                                   (mm_interconnect_0_cam_ctrl_slave_writedata),                 //                                                     .writedata
		.cam_ctrl_slave_chipselect                                  (mm_interconnect_0_cam_ctrl_slave_chipselect),                //                                                     .chipselect
		.i2c_ctrl_slave_address                                     (mm_interconnect_0_i2c_ctrl_slave_address),                   //                                       i2c_ctrl_slave.address
		.i2c_ctrl_slave_write                                       (mm_interconnect_0_i2c_ctrl_slave_write),                     //                                                     .write
		.i2c_ctrl_slave_readdata                                    (mm_interconnect_0_i2c_ctrl_slave_readdata),                  //                                                     .readdata
		.i2c_ctrl_slave_writedata                                   (mm_interconnect_0_i2c_ctrl_slave_writedata),                 //                                                     .writedata
		.i2c_ctrl_slave_byteenable                                  (mm_interconnect_0_i2c_ctrl_slave_byteenable),                //                                                     .byteenable
		.i2c_ctrl_slave_chipselect                                  (mm_interconnect_0_i2c_ctrl_slave_chipselect),                //                                                     .chipselect
		.jtag_uart_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //                          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                                     .write
		.jtag_uart_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                                     .read
		.jtag_uart_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                                     .chipselect
		.lcd_ctrl_slave_address                                     (mm_interconnect_0_lcd_ctrl_slave_address),                   //                                       lcd_ctrl_slave.address
		.lcd_ctrl_slave_write                                       (mm_interconnect_0_lcd_ctrl_slave_write),                     //                                                     .write
		.lcd_ctrl_slave_read                                        (mm_interconnect_0_lcd_ctrl_slave_read),                      //                                                     .read
		.lcd_ctrl_slave_readdata                                    (mm_interconnect_0_lcd_ctrl_slave_readdata),                  //                                                     .readdata
		.lcd_ctrl_slave_writedata                                   (mm_interconnect_0_lcd_ctrl_slave_writedata),                 //                                                     .writedata
		.lcd_ctrl_slave_waitrequest                                 (mm_interconnect_0_lcd_ctrl_slave_waitrequest),               //                                                     .waitrequest
		.lcd_ctrl_slave_chipselect                                  (mm_interconnect_0_lcd_ctrl_slave_chipselect),                //                                                     .chipselect
		.nios2_gen2_0_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //                         nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                                     .write
		.nios2_gen2_0_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                                     .read
		.nios2_gen2_0_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                                     .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                                     .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                                     .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                                     .debugaccess
		.pio_0_s1_address                                           (mm_interconnect_0_pio_0_s1_address),                         //                                             pio_0_s1.address
		.pio_0_s1_readdata                                          (mm_interconnect_0_pio_0_s1_readdata),                        //                                                     .readdata
		.ProfileTimer_s1_address                                    (mm_interconnect_0_profiletimer_s1_address),                  //                                      ProfileTimer_s1.address
		.ProfileTimer_s1_write                                      (mm_interconnect_0_profiletimer_s1_write),                    //                                                     .write
		.ProfileTimer_s1_readdata                                   (mm_interconnect_0_profiletimer_s1_readdata),                 //                                                     .readdata
		.ProfileTimer_s1_writedata                                  (mm_interconnect_0_profiletimer_s1_writedata),                //                                                     .writedata
		.ProfileTimer_s1_chipselect                                 (mm_interconnect_0_profiletimer_s1_chipselect),               //                                                     .chipselect
		.sdram_ctrl_s1_address                                      (mm_interconnect_0_sdram_ctrl_s1_address),                    //                                        sdram_ctrl_s1.address
		.sdram_ctrl_s1_write                                        (mm_interconnect_0_sdram_ctrl_s1_write),                      //                                                     .write
		.sdram_ctrl_s1_read                                         (mm_interconnect_0_sdram_ctrl_s1_read),                       //                                                     .read
		.sdram_ctrl_s1_readdata                                     (mm_interconnect_0_sdram_ctrl_s1_readdata),                   //                                                     .readdata
		.sdram_ctrl_s1_writedata                                    (mm_interconnect_0_sdram_ctrl_s1_writedata),                  //                                                     .writedata
		.sdram_ctrl_s1_byteenable                                   (mm_interconnect_0_sdram_ctrl_s1_byteenable),                 //                                                     .byteenable
		.sdram_ctrl_s1_readdatavalid                                (mm_interconnect_0_sdram_ctrl_s1_readdatavalid),              //                                                     .readdatavalid
		.sdram_ctrl_s1_waitrequest                                  (mm_interconnect_0_sdram_ctrl_s1_waitrequest),                //                                                     .waitrequest
		.sdram_ctrl_s1_chipselect                                   (mm_interconnect_0_sdram_ctrl_s1_chipselect),                 //                                                     .chipselect
		.sysid_control_slave_address                                (mm_interconnect_0_sysid_control_slave_address),              //                                  sysid_control_slave.address
		.sysid_control_slave_readdata                               (mm_interconnect_0_sysid_control_slave_readdata),             //                                                     .readdata
		.Systimer_s1_address                                        (mm_interconnect_0_systimer_s1_address),                      //                                          Systimer_s1.address
		.Systimer_s1_write                                          (mm_interconnect_0_systimer_s1_write),                        //                                                     .write
		.Systimer_s1_readdata                                       (mm_interconnect_0_systimer_s1_readdata),                     //                                                     .readdata
		.Systimer_s1_writedata                                      (mm_interconnect_0_systimer_s1_writedata),                    //                                                     .writedata
		.Systimer_s1_chipselect                                     (mm_interconnect_0_systimer_s1_chipselect),                   //                                                     .chipselect
		.vga_dma_0_slave_address                                    (mm_interconnect_0_vga_dma_0_slave_address),                  //                                      vga_dma_0_slave.address
		.vga_dma_0_slave_write                                      (mm_interconnect_0_vga_dma_0_slave_write),                    //                                                     .write
		.vga_dma_0_slave_writedata                                  (mm_interconnect_0_vga_dma_0_slave_writedata),                //                                                     .writedata
		.vga_dma_0_slave_chipselect                                 (mm_interconnect_0_vga_dma_0_slave_chipselect)                //                                                     .chipselect
	);

	base_system_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
